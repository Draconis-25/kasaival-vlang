module lyra

pub const (
	game_width  = 1920
	game_height = 1080
)
