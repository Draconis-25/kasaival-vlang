module plants
