module stages

fn desert_props() []Scene {
	mut one := Scene{}
	one.add_width = 20000
	one.color_scheme = [
	// water
	[80, 100, 60, 90, 140, 180],
	[100, 120, 80, 110, 140, 190],
	[100, 140, 90, 120, 160, 205],
	[130, 160, 120, 130, 160, 205],
	[140, 170, 120, 140, 140, 175],
	// shore
		[150, 180, 120, 140, 130, 155],
		[180, 200, 130, 150, 120, 135],
		// sand
		[190, 210, 140, 160, 100, 125],
		[190, 210, 140, 160, 100, 125],
		[190, 210, 140, 160, 100, 125],
		[200, 220, 150, 180, 80, 105],
		[200, 220, 150, 180, 80, 105],
		[200, 220, 150, 180, 80, 105],
		[200, 220, 150, 180, 80, 105],
	// desert
		[190, 200, 130, 150, 80, 105],
		[170, 200, 115, 140, 80, 84],
		[200, 220, 115, 140, 75, 80],
		[220, 230, 105, 122, 54, 80],
	// shore
	[220, 230, 105, 122, 74, 90],
	[200, 220, 115, 140, 85, 100],
	[170, 200, 115, 140, 100, 124],
	]
	return [one]
}
