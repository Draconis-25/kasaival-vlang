module plants

pub fn saguaro(mut self Core)  {
	self.cs_branch = [125, 178, 122, 160, 76, 90]
	self.cs_leaf = [150, 204, 190, 230, 159, 178]
	self.change_color = [-10, -25, -20]
	self.grow_time = 20
	self.max_row = 7
	self.w = 14
	self.h = 42
	self.split_chance = 40
}
