module stages

fn grassland() []Scene {
	mut scene := Scene{}
	scene.ground.width += 3000
	scene.ground.cs = [
		// grassland
		[80, 140, 100, 150, 40, 64],
		[80, 160, 135, 170, 55, 60],
	]
	// add saguaro spawner to spawners
	scene.spawners << get_spawner(.oak, 100)
	// add mob spawner

	// set Music
	scene.music = 'spring/map.ogg'

	// set background
	scene.background = 'grassland'
	// return all scenes
	return [scene]
}
